library verilog;
use verilog.vl_types.all;
entity Secador_vlg_check_tst is
    port(
        DATA_MISO       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Secador_vlg_check_tst;
