-- megafunction wizard: %ALTFP_COMPARE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altfp_compare 

-- ============================================================
-- File Name: altfp_compare_PWM_EN.vhd
-- Megafunction Name(s):
-- 			altfp_compare
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.0 Build 156 04/24/2013 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_compare CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" PIPELINE=1 WIDTH_EXP=8 WIDTH_MAN=23 agb clock dataa datab
--VERSION_BEGIN 13.0 cbx_altfp_compare 2013:04:24:18:05:29:SJ cbx_cycloneii 2013:04:24:18:05:30:SJ cbx_lpm_add_sub 2013:04:24:18:05:30:SJ cbx_lpm_compare 2013:04:24:18:05:30:SJ cbx_mgl 2013:04:24:18:40:34:SJ cbx_stratix 2013:04:24:18:05:30:SJ cbx_stratixii 2013:04:24:18:05:30:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_compare 4 reg 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_compare_PWM_EN_altfp_compare_h3b IS 
	 PORT 
	 ( 
		 agb	:	OUT  STD_LOGIC;
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END altfp_compare_PWM_EN_altfp_compare_h3b;

 ARCHITECTURE RTL OF altfp_compare_PWM_EN_altfp_compare_h3b IS

	 SIGNAL	 out_agb_w_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cmpr1_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr1_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr2_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr2_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr3_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr3_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr4_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr4_agb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w304w305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_agb_w_dffe2_wo314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_flip_outputs_dffe2_wo310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range11w17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range21w27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range31w37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range41w47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range51w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range61w67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range71w77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range14w19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range24w29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range34w39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range44w49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range54w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range64w69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range74w79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_aeb_range233w245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_aeb_range237w247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_aeb_range241w249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_eq_grp_range251w253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_eq_grp_range251w259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_eq_grp_range254w255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_eq_grp_range254w261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_eq_grp_range256w263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_both_inputs_zero_dffe2_wo312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_a_not_zero_dffe1_wo293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_agb_w_dffe2_wo309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_b_not_zero_dffe1_wo294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_dataa_zero_w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_datab_zero_w298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_out_aeb_w308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_out_unordered_w302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w304w305w306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range141w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range147w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range157w158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range163w164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range169w170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range175w176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range181w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range187w188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range193w194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range87w88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range199w200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range205w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range211w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range11w12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range21w22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range31w32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range41w42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range51w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range61w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range93w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range71w72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range99w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range105w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range111w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range117w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range123w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range129w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range135w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range144w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range150w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range160w161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range166w167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range172w173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range178w179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range184w185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range190w191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range196w197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range90w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range202w203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range208w209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range214w215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range14w15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range24w25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range34w35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range44w45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range54w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range64w65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range96w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range74w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range102w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range108w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range114w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range120w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range126w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range132w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range138w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_agb_tmp_w_range265w267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_agb_tmp_w_range268w269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_agb_tmp_w_range270w271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_not_zero_dffe1_wo_range285w286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_not_zero_dffe1_wo_range288w289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_adjusted_dffe2_wi :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_adjusted_dffe2_wo :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_adjusted_w :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_dffe1_wi :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_dffe1_wo :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_w :	STD_LOGIC;
	 SIGNAL  aligned_dataa_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  aligned_datab_sign_adjusted_dffe2_wi :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_adjusted_dffe2_wo :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_adjusted_w :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_dffe1_wi :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_dffe1_wo :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_w :	STD_LOGIC;
	 SIGNAL  aligned_datab_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  both_inputs_zero :	STD_LOGIC;
	 SIGNAL  both_inputs_zero_dffe2_wi :	STD_LOGIC;
	 SIGNAL  both_inputs_zero_dffe2_wo :	STD_LOGIC;
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  exp_a_all_one_dffe1_wi :	STD_LOGIC;
	 SIGNAL  exp_a_all_one_dffe1_wo :	STD_LOGIC;
	 SIGNAL  exp_a_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_a_not_zero_dffe1_wi :	STD_LOGIC;
	 SIGNAL  exp_a_not_zero_dffe1_wo :	STD_LOGIC;
	 SIGNAL  exp_a_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_aeb :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  exp_aeb_tmp_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  exp_aeb_w :	STD_LOGIC;
	 SIGNAL  exp_aeb_w_dffe2_wi :	STD_LOGIC;
	 SIGNAL  exp_aeb_w_dffe2_wo :	STD_LOGIC;
	 SIGNAL  exp_agb :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  exp_agb_tmp_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  exp_agb_w :	STD_LOGIC;
	 SIGNAL  exp_agb_w_dffe2_wi :	STD_LOGIC;
	 SIGNAL  exp_agb_w_dffe2_wo :	STD_LOGIC;
	 SIGNAL  exp_b_all_one_dffe1_wi :	STD_LOGIC;
	 SIGNAL  exp_b_all_one_dffe1_wo :	STD_LOGIC;
	 SIGNAL  exp_b_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_b_not_zero_dffe1_wi :	STD_LOGIC;
	 SIGNAL  exp_b_not_zero_dffe1_wo :	STD_LOGIC;
	 SIGNAL  exp_b_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_eq_grp :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  exp_eq_gt_grp :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  flip_outputs_dffe2_wi :	STD_LOGIC;
	 SIGNAL  flip_outputs_dffe2_wo :	STD_LOGIC;
	 SIGNAL  flip_outputs_w :	STD_LOGIC;
	 SIGNAL  input_dataa_nan_dffe2_wi :	STD_LOGIC;
	 SIGNAL  input_dataa_nan_dffe2_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_nan_w :	STD_LOGIC;
	 SIGNAL  input_dataa_zero_w :	STD_LOGIC;
	 SIGNAL  input_datab_nan_dffe2_wi :	STD_LOGIC;
	 SIGNAL  input_datab_nan_dffe2_wo :	STD_LOGIC;
	 SIGNAL  input_datab_nan_w :	STD_LOGIC;
	 SIGNAL  input_datab_zero_w :	STD_LOGIC;
	 SIGNAL  man_a_not_zero_dffe1_wi :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_a_not_zero_dffe1_wo :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_a_not_zero_merge_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_a_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_not_zero_dffe1_wi :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_b_not_zero_dffe1_wo :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_b_not_zero_merge_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_b_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  out_aeb_w :	STD_LOGIC;
	 SIGNAL  out_agb_dffe3_wi :	STD_LOGIC;
	 SIGNAL  out_agb_dffe3_wo :	STD_LOGIC;
	 SIGNAL  out_agb_w :	STD_LOGIC;
	 SIGNAL  out_unordered_w :	STD_LOGIC;
	 SIGNAL  wire_w_dataa_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_range233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_range237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_range241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_tmp_w_range243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_tmp_w_range246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_tmp_w_range248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_range234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_range238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_range242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_tmp_w_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_tmp_w_range268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_tmp_w_range270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_grp_range251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_grp_range254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_grp_range256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_gt_grp_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_gt_grp_range262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_gt_grp_range264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_dffe1_wo_range285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_merge_w_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_dffe1_wo_range288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_merge_w_range283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w304w305w(0) <= wire_w304w(0) AND exp_aeb_w_dffe2_wo;
	wire_w316w(0) <= wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo313w(0) AND aligned_datab_sign_adjusted_dffe2_wo;
	wire_w_lg_exp_agb_w_dffe2_wo314w(0) <= exp_agb_w_dffe2_wo AND wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo313w(0);
	wire_w_lg_flip_outputs_dffe2_wo310w(0) <= flip_outputs_dffe2_wo AND wire_w_lg_exp_agb_w_dffe2_wo309w(0);
	wire_w_lg_w_dataa_range11w17w(0) <= wire_w_dataa_range11w(0) AND wire_w_exp_a_all_one_w_range7w(0);
	wire_w_lg_w_dataa_range21w27w(0) <= wire_w_dataa_range21w(0) AND wire_w_exp_a_all_one_w_range18w(0);
	wire_w_lg_w_dataa_range31w37w(0) <= wire_w_dataa_range31w(0) AND wire_w_exp_a_all_one_w_range28w(0);
	wire_w_lg_w_dataa_range41w47w(0) <= wire_w_dataa_range41w(0) AND wire_w_exp_a_all_one_w_range38w(0);
	wire_w_lg_w_dataa_range51w57w(0) <= wire_w_dataa_range51w(0) AND wire_w_exp_a_all_one_w_range48w(0);
	wire_w_lg_w_dataa_range61w67w(0) <= wire_w_dataa_range61w(0) AND wire_w_exp_a_all_one_w_range58w(0);
	wire_w_lg_w_dataa_range71w77w(0) <= wire_w_dataa_range71w(0) AND wire_w_exp_a_all_one_w_range68w(0);
	wire_w_lg_w_datab_range14w19w(0) <= wire_w_datab_range14w(0) AND wire_w_exp_b_all_one_w_range9w(0);
	wire_w_lg_w_datab_range24w29w(0) <= wire_w_datab_range24w(0) AND wire_w_exp_b_all_one_w_range20w(0);
	wire_w_lg_w_datab_range34w39w(0) <= wire_w_datab_range34w(0) AND wire_w_exp_b_all_one_w_range30w(0);
	wire_w_lg_w_datab_range44w49w(0) <= wire_w_datab_range44w(0) AND wire_w_exp_b_all_one_w_range40w(0);
	wire_w_lg_w_datab_range54w59w(0) <= wire_w_datab_range54w(0) AND wire_w_exp_b_all_one_w_range50w(0);
	wire_w_lg_w_datab_range64w69w(0) <= wire_w_datab_range64w(0) AND wire_w_exp_b_all_one_w_range60w(0);
	wire_w_lg_w_datab_range74w79w(0) <= wire_w_datab_range74w(0) AND wire_w_exp_b_all_one_w_range70w(0);
	wire_w_lg_w_exp_aeb_range233w245w(0) <= wire_w_exp_aeb_range233w(0) AND wire_w_exp_aeb_tmp_w_range243w(0);
	wire_w_lg_w_exp_aeb_range237w247w(0) <= wire_w_exp_aeb_range237w(0) AND wire_w_exp_aeb_tmp_w_range246w(0);
	wire_w_lg_w_exp_aeb_range241w249w(0) <= wire_w_exp_aeb_range241w(0) AND wire_w_exp_aeb_tmp_w_range248w(0);
	wire_w_lg_w_exp_eq_grp_range251w253w(0) <= wire_w_exp_eq_grp_range251w(0) AND wire_w_exp_aeb_range233w(0);
	wire_w_lg_w_exp_eq_grp_range251w259w(0) <= wire_w_exp_eq_grp_range251w(0) AND wire_w_exp_agb_range234w(0);
	wire_w_lg_w_exp_eq_grp_range254w255w(0) <= wire_w_exp_eq_grp_range254w(0) AND wire_w_exp_aeb_range237w(0);
	wire_w_lg_w_exp_eq_grp_range254w261w(0) <= wire_w_exp_eq_grp_range254w(0) AND wire_w_exp_agb_range238w(0);
	wire_w_lg_w_exp_eq_grp_range256w263w(0) <= wire_w_exp_eq_grp_range256w(0) AND wire_w_exp_agb_range242w(0);
	wire_w304w(0) <= NOT wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo303w(0);
	wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo313w(0) <= NOT aligned_dataa_sign_adjusted_dffe2_wo;
	wire_w_lg_both_inputs_zero_dffe2_wo312w(0) <= NOT both_inputs_zero_dffe2_wo;
	wire_w_lg_exp_a_not_zero_dffe1_wo293w(0) <= NOT exp_a_not_zero_dffe1_wo;
	wire_w_lg_exp_agb_w_dffe2_wo309w(0) <= NOT exp_agb_w_dffe2_wo;
	wire_w_lg_exp_b_not_zero_dffe1_wo294w(0) <= NOT exp_b_not_zero_dffe1_wo;
	wire_w_lg_input_dataa_zero_w296w(0) <= NOT input_dataa_zero_w;
	wire_w_lg_input_datab_zero_w298w(0) <= NOT input_datab_zero_w;
	wire_w_lg_out_aeb_w308w(0) <= NOT out_aeb_w;
	wire_w_lg_out_unordered_w302w(0) <= NOT out_unordered_w;
	wire_w_lg_w_lg_w304w305w306w(0) <= wire_w_lg_w304w305w(0) OR both_inputs_zero_dffe2_wo;
	wire_w_lg_w_dataa_range141w142w(0) <= wire_w_dataa_range141w(0) OR wire_w_man_a_not_zero_w_range137w(0);
	wire_w_lg_w_dataa_range147w148w(0) <= wire_w_dataa_range147w(0) OR wire_w_man_a_not_zero_w_range143w(0);
	wire_w_lg_w_dataa_range157w158w(0) <= wire_w_dataa_range157w(0) OR wire_w_man_a_not_zero_w_range154w(0);
	wire_w_lg_w_dataa_range163w164w(0) <= wire_w_dataa_range163w(0) OR wire_w_man_a_not_zero_w_range159w(0);
	wire_w_lg_w_dataa_range169w170w(0) <= wire_w_dataa_range169w(0) OR wire_w_man_a_not_zero_w_range165w(0);
	wire_w_lg_w_dataa_range175w176w(0) <= wire_w_dataa_range175w(0) OR wire_w_man_a_not_zero_w_range171w(0);
	wire_w_lg_w_dataa_range181w182w(0) <= wire_w_dataa_range181w(0) OR wire_w_man_a_not_zero_w_range177w(0);
	wire_w_lg_w_dataa_range187w188w(0) <= wire_w_dataa_range187w(0) OR wire_w_man_a_not_zero_w_range183w(0);
	wire_w_lg_w_dataa_range193w194w(0) <= wire_w_dataa_range193w(0) OR wire_w_man_a_not_zero_w_range189w(0);
	wire_w_lg_w_dataa_range87w88w(0) <= wire_w_dataa_range87w(0) OR wire_w_man_a_not_zero_w_range82w(0);
	wire_w_lg_w_dataa_range199w200w(0) <= wire_w_dataa_range199w(0) OR wire_w_man_a_not_zero_w_range195w(0);
	wire_w_lg_w_dataa_range205w206w(0) <= wire_w_dataa_range205w(0) OR wire_w_man_a_not_zero_w_range201w(0);
	wire_w_lg_w_dataa_range211w212w(0) <= wire_w_dataa_range211w(0) OR wire_w_man_a_not_zero_w_range207w(0);
	wire_w_lg_w_dataa_range11w12w(0) <= wire_w_dataa_range11w(0) OR wire_w_exp_a_not_zero_w_range2w(0);
	wire_w_lg_w_dataa_range21w22w(0) <= wire_w_dataa_range21w(0) OR wire_w_exp_a_not_zero_w_range13w(0);
	wire_w_lg_w_dataa_range31w32w(0) <= wire_w_dataa_range31w(0) OR wire_w_exp_a_not_zero_w_range23w(0);
	wire_w_lg_w_dataa_range41w42w(0) <= wire_w_dataa_range41w(0) OR wire_w_exp_a_not_zero_w_range33w(0);
	wire_w_lg_w_dataa_range51w52w(0) <= wire_w_dataa_range51w(0) OR wire_w_exp_a_not_zero_w_range43w(0);
	wire_w_lg_w_dataa_range61w62w(0) <= wire_w_dataa_range61w(0) OR wire_w_exp_a_not_zero_w_range53w(0);
	wire_w_lg_w_dataa_range93w94w(0) <= wire_w_dataa_range93w(0) OR wire_w_man_a_not_zero_w_range89w(0);
	wire_w_lg_w_dataa_range71w72w(0) <= wire_w_dataa_range71w(0) OR wire_w_exp_a_not_zero_w_range63w(0);
	wire_w_lg_w_dataa_range99w100w(0) <= wire_w_dataa_range99w(0) OR wire_w_man_a_not_zero_w_range95w(0);
	wire_w_lg_w_dataa_range105w106w(0) <= wire_w_dataa_range105w(0) OR wire_w_man_a_not_zero_w_range101w(0);
	wire_w_lg_w_dataa_range111w112w(0) <= wire_w_dataa_range111w(0) OR wire_w_man_a_not_zero_w_range107w(0);
	wire_w_lg_w_dataa_range117w118w(0) <= wire_w_dataa_range117w(0) OR wire_w_man_a_not_zero_w_range113w(0);
	wire_w_lg_w_dataa_range123w124w(0) <= wire_w_dataa_range123w(0) OR wire_w_man_a_not_zero_w_range119w(0);
	wire_w_lg_w_dataa_range129w130w(0) <= wire_w_dataa_range129w(0) OR wire_w_man_a_not_zero_w_range125w(0);
	wire_w_lg_w_dataa_range135w136w(0) <= wire_w_dataa_range135w(0) OR wire_w_man_a_not_zero_w_range131w(0);
	wire_w_lg_w_datab_range144w145w(0) <= wire_w_datab_range144w(0) OR wire_w_man_b_not_zero_w_range140w(0);
	wire_w_lg_w_datab_range150w151w(0) <= wire_w_datab_range150w(0) OR wire_w_man_b_not_zero_w_range146w(0);
	wire_w_lg_w_datab_range160w161w(0) <= wire_w_datab_range160w(0) OR wire_w_man_b_not_zero_w_range156w(0);
	wire_w_lg_w_datab_range166w167w(0) <= wire_w_datab_range166w(0) OR wire_w_man_b_not_zero_w_range162w(0);
	wire_w_lg_w_datab_range172w173w(0) <= wire_w_datab_range172w(0) OR wire_w_man_b_not_zero_w_range168w(0);
	wire_w_lg_w_datab_range178w179w(0) <= wire_w_datab_range178w(0) OR wire_w_man_b_not_zero_w_range174w(0);
	wire_w_lg_w_datab_range184w185w(0) <= wire_w_datab_range184w(0) OR wire_w_man_b_not_zero_w_range180w(0);
	wire_w_lg_w_datab_range190w191w(0) <= wire_w_datab_range190w(0) OR wire_w_man_b_not_zero_w_range186w(0);
	wire_w_lg_w_datab_range196w197w(0) <= wire_w_datab_range196w(0) OR wire_w_man_b_not_zero_w_range192w(0);
	wire_w_lg_w_datab_range90w91w(0) <= wire_w_datab_range90w(0) OR wire_w_man_b_not_zero_w_range85w(0);
	wire_w_lg_w_datab_range202w203w(0) <= wire_w_datab_range202w(0) OR wire_w_man_b_not_zero_w_range198w(0);
	wire_w_lg_w_datab_range208w209w(0) <= wire_w_datab_range208w(0) OR wire_w_man_b_not_zero_w_range204w(0);
	wire_w_lg_w_datab_range214w215w(0) <= wire_w_datab_range214w(0) OR wire_w_man_b_not_zero_w_range210w(0);
	wire_w_lg_w_datab_range14w15w(0) <= wire_w_datab_range14w(0) OR wire_w_exp_b_not_zero_w_range5w(0);
	wire_w_lg_w_datab_range24w25w(0) <= wire_w_datab_range24w(0) OR wire_w_exp_b_not_zero_w_range16w(0);
	wire_w_lg_w_datab_range34w35w(0) <= wire_w_datab_range34w(0) OR wire_w_exp_b_not_zero_w_range26w(0);
	wire_w_lg_w_datab_range44w45w(0) <= wire_w_datab_range44w(0) OR wire_w_exp_b_not_zero_w_range36w(0);
	wire_w_lg_w_datab_range54w55w(0) <= wire_w_datab_range54w(0) OR wire_w_exp_b_not_zero_w_range46w(0);
	wire_w_lg_w_datab_range64w65w(0) <= wire_w_datab_range64w(0) OR wire_w_exp_b_not_zero_w_range56w(0);
	wire_w_lg_w_datab_range96w97w(0) <= wire_w_datab_range96w(0) OR wire_w_man_b_not_zero_w_range92w(0);
	wire_w_lg_w_datab_range74w75w(0) <= wire_w_datab_range74w(0) OR wire_w_exp_b_not_zero_w_range66w(0);
	wire_w_lg_w_datab_range102w103w(0) <= wire_w_datab_range102w(0) OR wire_w_man_b_not_zero_w_range98w(0);
	wire_w_lg_w_datab_range108w109w(0) <= wire_w_datab_range108w(0) OR wire_w_man_b_not_zero_w_range104w(0);
	wire_w_lg_w_datab_range114w115w(0) <= wire_w_datab_range114w(0) OR wire_w_man_b_not_zero_w_range110w(0);
	wire_w_lg_w_datab_range120w121w(0) <= wire_w_datab_range120w(0) OR wire_w_man_b_not_zero_w_range116w(0);
	wire_w_lg_w_datab_range126w127w(0) <= wire_w_datab_range126w(0) OR wire_w_man_b_not_zero_w_range122w(0);
	wire_w_lg_w_datab_range132w133w(0) <= wire_w_datab_range132w(0) OR wire_w_man_b_not_zero_w_range128w(0);
	wire_w_lg_w_datab_range138w139w(0) <= wire_w_datab_range138w(0) OR wire_w_man_b_not_zero_w_range134w(0);
	wire_w_lg_w_exp_agb_tmp_w_range265w267w(0) <= wire_w_exp_agb_tmp_w_range265w(0) OR wire_w_exp_eq_gt_grp_range260w(0);
	wire_w_lg_w_exp_agb_tmp_w_range268w269w(0) <= wire_w_exp_agb_tmp_w_range268w(0) OR wire_w_exp_eq_gt_grp_range262w(0);
	wire_w_lg_w_exp_agb_tmp_w_range270w271w(0) <= wire_w_exp_agb_tmp_w_range270w(0) OR wire_w_exp_eq_gt_grp_range264w(0);
	wire_w_lg_w_man_a_not_zero_dffe1_wo_range285w286w(0) <= wire_w_man_a_not_zero_dffe1_wo_range285w(0) OR wire_w_man_a_not_zero_merge_w_range280w(0);
	wire_w_lg_w_man_b_not_zero_dffe1_wo_range288w289w(0) <= wire_w_man_b_not_zero_dffe1_wo_range288w(0) OR wire_w_man_b_not_zero_merge_w_range283w(0);
	wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo303w(0) <= aligned_dataa_sign_adjusted_dffe2_wo XOR aligned_datab_sign_adjusted_dffe2_wo;
	aclr <= '0';
	agb <= out_agb_dffe3_wo;
	aligned_dataa_sign_adjusted_dffe2_wi <= aligned_dataa_sign_adjusted_w;
	aligned_dataa_sign_adjusted_dffe2_wo <= aligned_dataa_sign_adjusted_dffe2_wi;
	aligned_dataa_sign_adjusted_w <= (aligned_dataa_sign_dffe1_wo AND wire_w_lg_input_dataa_zero_w296w(0));
	aligned_dataa_sign_dffe1_wi <= aligned_dataa_sign_w;
	aligned_dataa_sign_dffe1_wo <= aligned_dataa_sign_dffe1_wi;
	aligned_dataa_sign_w <= dataa(31);
	aligned_dataa_w <= ( dataa(30 DOWNTO 0));
	aligned_datab_sign_adjusted_dffe2_wi <= aligned_datab_sign_adjusted_w;
	aligned_datab_sign_adjusted_dffe2_wo <= aligned_datab_sign_adjusted_dffe2_wi;
	aligned_datab_sign_adjusted_w <= (aligned_datab_sign_dffe1_wo AND wire_w_lg_input_datab_zero_w298w(0));
	aligned_datab_sign_dffe1_wi <= aligned_datab_sign_w;
	aligned_datab_sign_dffe1_wo <= aligned_datab_sign_dffe1_wi;
	aligned_datab_sign_w <= datab(31);
	aligned_datab_w <= ( datab(30 DOWNTO 0));
	both_inputs_zero <= (input_dataa_zero_w AND input_datab_zero_w);
	both_inputs_zero_dffe2_wi <= both_inputs_zero;
	both_inputs_zero_dffe2_wo <= both_inputs_zero_dffe2_wi;
	clk_en <= '1';
	exp_a_all_one_dffe1_wi <= exp_a_all_one_w(7);
	exp_a_all_one_dffe1_wo <= exp_a_all_one_dffe1_wi;
	exp_a_all_one_w <= ( wire_w_lg_w_dataa_range71w77w & wire_w_lg_w_dataa_range61w67w & wire_w_lg_w_dataa_range51w57w & wire_w_lg_w_dataa_range41w47w & wire_w_lg_w_dataa_range31w37w & wire_w_lg_w_dataa_range21w27w & wire_w_lg_w_dataa_range11w17w & dataa(23));
	exp_a_not_zero_dffe1_wi <= exp_a_not_zero_w(7);
	exp_a_not_zero_dffe1_wo <= exp_a_not_zero_dffe1_wi;
	exp_a_not_zero_w <= ( wire_w_lg_w_dataa_range71w72w & wire_w_lg_w_dataa_range61w62w & wire_w_lg_w_dataa_range51w52w & wire_w_lg_w_dataa_range41w42w & wire_w_lg_w_dataa_range31w32w & wire_w_lg_w_dataa_range21w22w & wire_w_lg_w_dataa_range11w12w & dataa(23));
	exp_aeb <= ( wire_cmpr4_aeb & wire_cmpr3_aeb & wire_cmpr2_aeb & wire_cmpr1_aeb);
	exp_aeb_tmp_w <= ( wire_w_lg_w_exp_aeb_range241w249w & wire_w_lg_w_exp_aeb_range237w247w & wire_w_lg_w_exp_aeb_range233w245w & exp_aeb(0));
	exp_aeb_w <= exp_aeb_tmp_w(3);
	exp_aeb_w_dffe2_wi <= exp_aeb_w;
	exp_aeb_w_dffe2_wo <= exp_aeb_w_dffe2_wi;
	exp_agb <= ( wire_cmpr4_agb & wire_cmpr3_agb & wire_cmpr2_agb & wire_cmpr1_agb);
	exp_agb_tmp_w <= ( wire_w_lg_w_exp_agb_tmp_w_range270w271w & wire_w_lg_w_exp_agb_tmp_w_range268w269w & wire_w_lg_w_exp_agb_tmp_w_range265w267w & exp_eq_gt_grp(0));
	exp_agb_w <= exp_agb_tmp_w(3);
	exp_agb_w_dffe2_wi <= exp_agb_w;
	exp_agb_w_dffe2_wo <= exp_agb_w_dffe2_wi;
	exp_b_all_one_dffe1_wi <= exp_b_all_one_w(7);
	exp_b_all_one_dffe1_wo <= exp_b_all_one_dffe1_wi;
	exp_b_all_one_w <= ( wire_w_lg_w_datab_range74w79w & wire_w_lg_w_datab_range64w69w & wire_w_lg_w_datab_range54w59w & wire_w_lg_w_datab_range44w49w & wire_w_lg_w_datab_range34w39w & wire_w_lg_w_datab_range24w29w & wire_w_lg_w_datab_range14w19w & datab(23));
	exp_b_not_zero_dffe1_wi <= exp_b_not_zero_w(7);
	exp_b_not_zero_dffe1_wo <= exp_b_not_zero_dffe1_wi;
	exp_b_not_zero_w <= ( wire_w_lg_w_datab_range74w75w & wire_w_lg_w_datab_range64w65w & wire_w_lg_w_datab_range54w55w & wire_w_lg_w_datab_range44w45w & wire_w_lg_w_datab_range34w35w & wire_w_lg_w_datab_range24w25w & wire_w_lg_w_datab_range14w15w & datab(23));
	exp_eq_grp <= ( wire_w_lg_w_exp_eq_grp_range254w255w & wire_w_lg_w_exp_eq_grp_range251w253w & exp_aeb(0));
	exp_eq_gt_grp <= ( wire_w_lg_w_exp_eq_grp_range256w263w & wire_w_lg_w_exp_eq_grp_range254w261w & wire_w_lg_w_exp_eq_grp_range251w259w & exp_agb(0));
	flip_outputs_dffe2_wi <= flip_outputs_w;
	flip_outputs_dffe2_wo <= flip_outputs_dffe2_wi;
	flip_outputs_w <= (aligned_dataa_sign_adjusted_w AND aligned_datab_sign_adjusted_w);
	input_dataa_nan_dffe2_wi <= input_dataa_nan_w;
	input_dataa_nan_dffe2_wo <= input_dataa_nan_dffe2_wi;
	input_dataa_nan_w <= (exp_a_all_one_dffe1_wo AND man_a_not_zero_merge_w(1));
	input_dataa_zero_w <= wire_w_lg_exp_a_not_zero_dffe1_wo293w(0);
	input_datab_nan_dffe2_wi <= input_datab_nan_w;
	input_datab_nan_dffe2_wo <= input_datab_nan_dffe2_wi;
	input_datab_nan_w <= (exp_b_all_one_dffe1_wo AND man_b_not_zero_merge_w(1));
	input_datab_zero_w <= wire_w_lg_exp_b_not_zero_dffe1_wo294w(0);
	man_a_not_zero_dffe1_wi <= ( man_a_not_zero_w(22) & man_a_not_zero_w(11));
	man_a_not_zero_dffe1_wo <= man_a_not_zero_dffe1_wi;
	man_a_not_zero_merge_w <= ( wire_w_lg_w_man_a_not_zero_dffe1_wo_range285w286w & man_a_not_zero_dffe1_wo(0));
	man_a_not_zero_w <= ( wire_w_lg_w_dataa_range211w212w & wire_w_lg_w_dataa_range205w206w & wire_w_lg_w_dataa_range199w200w & wire_w_lg_w_dataa_range193w194w & wire_w_lg_w_dataa_range187w188w & wire_w_lg_w_dataa_range181w182w & wire_w_lg_w_dataa_range175w176w & wire_w_lg_w_dataa_range169w170w & wire_w_lg_w_dataa_range163w164w & wire_w_lg_w_dataa_range157w158w & dataa(12) & wire_w_lg_w_dataa_range147w148w & wire_w_lg_w_dataa_range141w142w & wire_w_lg_w_dataa_range135w136w & wire_w_lg_w_dataa_range129w130w & wire_w_lg_w_dataa_range123w124w & wire_w_lg_w_dataa_range117w118w & wire_w_lg_w_dataa_range111w112w & wire_w_lg_w_dataa_range105w106w & wire_w_lg_w_dataa_range99w100w & wire_w_lg_w_dataa_range93w94w & wire_w_lg_w_dataa_range87w88w & dataa(0));
	man_b_not_zero_dffe1_wi <= ( man_b_not_zero_w(22) & man_b_not_zero_w(11));
	man_b_not_zero_dffe1_wo <= man_b_not_zero_dffe1_wi;
	man_b_not_zero_merge_w <= ( wire_w_lg_w_man_b_not_zero_dffe1_wo_range288w289w & man_b_not_zero_dffe1_wo(0));
	man_b_not_zero_w <= ( wire_w_lg_w_datab_range214w215w & wire_w_lg_w_datab_range208w209w & wire_w_lg_w_datab_range202w203w & wire_w_lg_w_datab_range196w197w & wire_w_lg_w_datab_range190w191w & wire_w_lg_w_datab_range184w185w & wire_w_lg_w_datab_range178w179w & wire_w_lg_w_datab_range172w173w & wire_w_lg_w_datab_range166w167w & wire_w_lg_w_datab_range160w161w & datab(12) & wire_w_lg_w_datab_range150w151w & wire_w_lg_w_datab_range144w145w & wire_w_lg_w_datab_range138w139w & wire_w_lg_w_datab_range132w133w & wire_w_lg_w_datab_range126w127w & wire_w_lg_w_datab_range120w121w & wire_w_lg_w_datab_range114w115w & wire_w_lg_w_datab_range108w109w & wire_w_lg_w_datab_range102w103w & wire_w_lg_w_datab_range96w97w & wire_w_lg_w_datab_range90w91w & datab(0));
	out_aeb_w <= (wire_w_lg_w_lg_w304w305w306w(0) AND wire_w_lg_out_unordered_w302w(0));
	out_agb_dffe3_wi <= out_agb_w;
	out_agb_dffe3_wo <= out_agb_w_dffe3;
	out_agb_w <= (((wire_w316w(0) OR (wire_w_lg_exp_agb_w_dffe2_wo314w(0) AND wire_w_lg_both_inputs_zero_dffe2_wo312w(0))) OR (wire_w_lg_flip_outputs_dffe2_wo310w(0) AND wire_w_lg_out_aeb_w308w(0))) AND wire_w_lg_out_unordered_w302w(0));
	out_unordered_w <= (input_dataa_nan_dffe2_wo OR input_datab_nan_dffe2_wo);
	wire_w_dataa_range141w(0) <= dataa(10);
	wire_w_dataa_range147w(0) <= dataa(11);
	wire_w_dataa_range157w(0) <= dataa(13);
	wire_w_dataa_range163w(0) <= dataa(14);
	wire_w_dataa_range169w(0) <= dataa(15);
	wire_w_dataa_range175w(0) <= dataa(16);
	wire_w_dataa_range181w(0) <= dataa(17);
	wire_w_dataa_range187w(0) <= dataa(18);
	wire_w_dataa_range193w(0) <= dataa(19);
	wire_w_dataa_range87w(0) <= dataa(1);
	wire_w_dataa_range199w(0) <= dataa(20);
	wire_w_dataa_range205w(0) <= dataa(21);
	wire_w_dataa_range211w(0) <= dataa(22);
	wire_w_dataa_range11w(0) <= dataa(24);
	wire_w_dataa_range21w(0) <= dataa(25);
	wire_w_dataa_range31w(0) <= dataa(26);
	wire_w_dataa_range41w(0) <= dataa(27);
	wire_w_dataa_range51w(0) <= dataa(28);
	wire_w_dataa_range61w(0) <= dataa(29);
	wire_w_dataa_range93w(0) <= dataa(2);
	wire_w_dataa_range71w(0) <= dataa(30);
	wire_w_dataa_range99w(0) <= dataa(3);
	wire_w_dataa_range105w(0) <= dataa(4);
	wire_w_dataa_range111w(0) <= dataa(5);
	wire_w_dataa_range117w(0) <= dataa(6);
	wire_w_dataa_range123w(0) <= dataa(7);
	wire_w_dataa_range129w(0) <= dataa(8);
	wire_w_dataa_range135w(0) <= dataa(9);
	wire_w_datab_range144w(0) <= datab(10);
	wire_w_datab_range150w(0) <= datab(11);
	wire_w_datab_range160w(0) <= datab(13);
	wire_w_datab_range166w(0) <= datab(14);
	wire_w_datab_range172w(0) <= datab(15);
	wire_w_datab_range178w(0) <= datab(16);
	wire_w_datab_range184w(0) <= datab(17);
	wire_w_datab_range190w(0) <= datab(18);
	wire_w_datab_range196w(0) <= datab(19);
	wire_w_datab_range90w(0) <= datab(1);
	wire_w_datab_range202w(0) <= datab(20);
	wire_w_datab_range208w(0) <= datab(21);
	wire_w_datab_range214w(0) <= datab(22);
	wire_w_datab_range14w(0) <= datab(24);
	wire_w_datab_range24w(0) <= datab(25);
	wire_w_datab_range34w(0) <= datab(26);
	wire_w_datab_range44w(0) <= datab(27);
	wire_w_datab_range54w(0) <= datab(28);
	wire_w_datab_range64w(0) <= datab(29);
	wire_w_datab_range96w(0) <= datab(2);
	wire_w_datab_range74w(0) <= datab(30);
	wire_w_datab_range102w(0) <= datab(3);
	wire_w_datab_range108w(0) <= datab(4);
	wire_w_datab_range114w(0) <= datab(5);
	wire_w_datab_range120w(0) <= datab(6);
	wire_w_datab_range126w(0) <= datab(7);
	wire_w_datab_range132w(0) <= datab(8);
	wire_w_datab_range138w(0) <= datab(9);
	wire_w_exp_a_all_one_w_range7w(0) <= exp_a_all_one_w(0);
	wire_w_exp_a_all_one_w_range18w(0) <= exp_a_all_one_w(1);
	wire_w_exp_a_all_one_w_range28w(0) <= exp_a_all_one_w(2);
	wire_w_exp_a_all_one_w_range38w(0) <= exp_a_all_one_w(3);
	wire_w_exp_a_all_one_w_range48w(0) <= exp_a_all_one_w(4);
	wire_w_exp_a_all_one_w_range58w(0) <= exp_a_all_one_w(5);
	wire_w_exp_a_all_one_w_range68w(0) <= exp_a_all_one_w(6);
	wire_w_exp_a_not_zero_w_range2w(0) <= exp_a_not_zero_w(0);
	wire_w_exp_a_not_zero_w_range13w(0) <= exp_a_not_zero_w(1);
	wire_w_exp_a_not_zero_w_range23w(0) <= exp_a_not_zero_w(2);
	wire_w_exp_a_not_zero_w_range33w(0) <= exp_a_not_zero_w(3);
	wire_w_exp_a_not_zero_w_range43w(0) <= exp_a_not_zero_w(4);
	wire_w_exp_a_not_zero_w_range53w(0) <= exp_a_not_zero_w(5);
	wire_w_exp_a_not_zero_w_range63w(0) <= exp_a_not_zero_w(6);
	wire_w_exp_aeb_range233w(0) <= exp_aeb(1);
	wire_w_exp_aeb_range237w(0) <= exp_aeb(2);
	wire_w_exp_aeb_range241w(0) <= exp_aeb(3);
	wire_w_exp_aeb_tmp_w_range243w(0) <= exp_aeb_tmp_w(0);
	wire_w_exp_aeb_tmp_w_range246w(0) <= exp_aeb_tmp_w(1);
	wire_w_exp_aeb_tmp_w_range248w(0) <= exp_aeb_tmp_w(2);
	wire_w_exp_agb_range234w(0) <= exp_agb(1);
	wire_w_exp_agb_range238w(0) <= exp_agb(2);
	wire_w_exp_agb_range242w(0) <= exp_agb(3);
	wire_w_exp_agb_tmp_w_range265w(0) <= exp_agb_tmp_w(0);
	wire_w_exp_agb_tmp_w_range268w(0) <= exp_agb_tmp_w(1);
	wire_w_exp_agb_tmp_w_range270w(0) <= exp_agb_tmp_w(2);
	wire_w_exp_b_all_one_w_range9w(0) <= exp_b_all_one_w(0);
	wire_w_exp_b_all_one_w_range20w(0) <= exp_b_all_one_w(1);
	wire_w_exp_b_all_one_w_range30w(0) <= exp_b_all_one_w(2);
	wire_w_exp_b_all_one_w_range40w(0) <= exp_b_all_one_w(3);
	wire_w_exp_b_all_one_w_range50w(0) <= exp_b_all_one_w(4);
	wire_w_exp_b_all_one_w_range60w(0) <= exp_b_all_one_w(5);
	wire_w_exp_b_all_one_w_range70w(0) <= exp_b_all_one_w(6);
	wire_w_exp_b_not_zero_w_range5w(0) <= exp_b_not_zero_w(0);
	wire_w_exp_b_not_zero_w_range16w(0) <= exp_b_not_zero_w(1);
	wire_w_exp_b_not_zero_w_range26w(0) <= exp_b_not_zero_w(2);
	wire_w_exp_b_not_zero_w_range36w(0) <= exp_b_not_zero_w(3);
	wire_w_exp_b_not_zero_w_range46w(0) <= exp_b_not_zero_w(4);
	wire_w_exp_b_not_zero_w_range56w(0) <= exp_b_not_zero_w(5);
	wire_w_exp_b_not_zero_w_range66w(0) <= exp_b_not_zero_w(6);
	wire_w_exp_eq_grp_range251w(0) <= exp_eq_grp(0);
	wire_w_exp_eq_grp_range254w(0) <= exp_eq_grp(1);
	wire_w_exp_eq_grp_range256w(0) <= exp_eq_grp(2);
	wire_w_exp_eq_gt_grp_range260w(0) <= exp_eq_gt_grp(1);
	wire_w_exp_eq_gt_grp_range262w(0) <= exp_eq_gt_grp(2);
	wire_w_exp_eq_gt_grp_range264w(0) <= exp_eq_gt_grp(3);
	wire_w_man_a_not_zero_dffe1_wo_range285w(0) <= man_a_not_zero_dffe1_wo(1);
	wire_w_man_a_not_zero_merge_w_range280w(0) <= man_a_not_zero_merge_w(0);
	wire_w_man_a_not_zero_w_range82w(0) <= man_a_not_zero_w(0);
	wire_w_man_a_not_zero_w_range143w(0) <= man_a_not_zero_w(10);
	wire_w_man_a_not_zero_w_range154w(0) <= man_a_not_zero_w(12);
	wire_w_man_a_not_zero_w_range159w(0) <= man_a_not_zero_w(13);
	wire_w_man_a_not_zero_w_range165w(0) <= man_a_not_zero_w(14);
	wire_w_man_a_not_zero_w_range171w(0) <= man_a_not_zero_w(15);
	wire_w_man_a_not_zero_w_range177w(0) <= man_a_not_zero_w(16);
	wire_w_man_a_not_zero_w_range183w(0) <= man_a_not_zero_w(17);
	wire_w_man_a_not_zero_w_range189w(0) <= man_a_not_zero_w(18);
	wire_w_man_a_not_zero_w_range195w(0) <= man_a_not_zero_w(19);
	wire_w_man_a_not_zero_w_range89w(0) <= man_a_not_zero_w(1);
	wire_w_man_a_not_zero_w_range201w(0) <= man_a_not_zero_w(20);
	wire_w_man_a_not_zero_w_range207w(0) <= man_a_not_zero_w(21);
	wire_w_man_a_not_zero_w_range95w(0) <= man_a_not_zero_w(2);
	wire_w_man_a_not_zero_w_range101w(0) <= man_a_not_zero_w(3);
	wire_w_man_a_not_zero_w_range107w(0) <= man_a_not_zero_w(4);
	wire_w_man_a_not_zero_w_range113w(0) <= man_a_not_zero_w(5);
	wire_w_man_a_not_zero_w_range119w(0) <= man_a_not_zero_w(6);
	wire_w_man_a_not_zero_w_range125w(0) <= man_a_not_zero_w(7);
	wire_w_man_a_not_zero_w_range131w(0) <= man_a_not_zero_w(8);
	wire_w_man_a_not_zero_w_range137w(0) <= man_a_not_zero_w(9);
	wire_w_man_b_not_zero_dffe1_wo_range288w(0) <= man_b_not_zero_dffe1_wo(1);
	wire_w_man_b_not_zero_merge_w_range283w(0) <= man_b_not_zero_merge_w(0);
	wire_w_man_b_not_zero_w_range85w(0) <= man_b_not_zero_w(0);
	wire_w_man_b_not_zero_w_range146w(0) <= man_b_not_zero_w(10);
	wire_w_man_b_not_zero_w_range156w(0) <= man_b_not_zero_w(12);
	wire_w_man_b_not_zero_w_range162w(0) <= man_b_not_zero_w(13);
	wire_w_man_b_not_zero_w_range168w(0) <= man_b_not_zero_w(14);
	wire_w_man_b_not_zero_w_range174w(0) <= man_b_not_zero_w(15);
	wire_w_man_b_not_zero_w_range180w(0) <= man_b_not_zero_w(16);
	wire_w_man_b_not_zero_w_range186w(0) <= man_b_not_zero_w(17);
	wire_w_man_b_not_zero_w_range192w(0) <= man_b_not_zero_w(18);
	wire_w_man_b_not_zero_w_range198w(0) <= man_b_not_zero_w(19);
	wire_w_man_b_not_zero_w_range92w(0) <= man_b_not_zero_w(1);
	wire_w_man_b_not_zero_w_range204w(0) <= man_b_not_zero_w(20);
	wire_w_man_b_not_zero_w_range210w(0) <= man_b_not_zero_w(21);
	wire_w_man_b_not_zero_w_range98w(0) <= man_b_not_zero_w(2);
	wire_w_man_b_not_zero_w_range104w(0) <= man_b_not_zero_w(3);
	wire_w_man_b_not_zero_w_range110w(0) <= man_b_not_zero_w(4);
	wire_w_man_b_not_zero_w_range116w(0) <= man_b_not_zero_w(5);
	wire_w_man_b_not_zero_w_range122w(0) <= man_b_not_zero_w(6);
	wire_w_man_b_not_zero_w_range128w(0) <= man_b_not_zero_w(7);
	wire_w_man_b_not_zero_w_range134w(0) <= man_b_not_zero_w(8);
	wire_w_man_b_not_zero_w_range140w(0) <= man_b_not_zero_w(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN out_agb_w_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN out_agb_w_dffe3 <= out_agb_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	cmpr1 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_cmpr1_aeb,
		agb => wire_cmpr1_agb,
		dataa => aligned_dataa_w(30 DOWNTO 23),
		datab => aligned_datab_w(30 DOWNTO 23)
	  );
	cmpr2 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_cmpr2_aeb,
		agb => wire_cmpr2_agb,
		dataa => aligned_dataa_w(22 DOWNTO 15),
		datab => aligned_datab_w(22 DOWNTO 15)
	  );
	cmpr3 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_cmpr3_aeb,
		agb => wire_cmpr3_agb,
		dataa => aligned_dataa_w(14 DOWNTO 7),
		datab => aligned_datab_w(14 DOWNTO 7)
	  );
	cmpr4 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 7
	  )
	  PORT MAP ( 
		aeb => wire_cmpr4_aeb,
		agb => wire_cmpr4_agb,
		dataa => aligned_dataa_w(6 DOWNTO 0),
		datab => aligned_datab_w(6 DOWNTO 0)
	  );

 END RTL; --altfp_compare_PWM_EN_altfp_compare_h3b
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altfp_compare_PWM_EN IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		agb		: OUT STD_LOGIC 
	);
END altfp_compare_PWM_EN;


ARCHITECTURE RTL OF altfp_compare_pwm_en IS

	SIGNAL sub_wire0	: STD_LOGIC ;



	COMPONENT altfp_compare_PWM_EN_altfp_compare_h3b
	PORT (
			agb	: OUT STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	agb    <= sub_wire0;

	altfp_compare_PWM_EN_altfp_compare_h3b_component : altfp_compare_PWM_EN_altfp_compare_h3b
	PORT MAP (
		clock => clock,
		dataa => dataa,
		datab => datab,
		agb => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: FPM_FORMAT NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "1"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: agb 0 0 0 0 OUTPUT NODEFVAL "agb"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: USED_PORT: datab 0 0 32 0 INPUT NODEFVAL "datab[31..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: CONNECT: @datab 0 0 32 0 datab 0 0 32 0
-- Retrieval info: CONNECT: agb 0 0 0 0 @agb 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_compare_PWM_EN.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_compare_PWM_EN.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_compare_PWM_EN.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_compare_PWM_EN.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_compare_PWM_EN_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
