-- megafunction wizard: %ALTFP_CONVERT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_CONVERT 

-- ============================================================
-- File Name: altfp_convert_INT_TO_FP.vhd
-- Megafunction Name(s):
-- 			ALTFP_CONVERT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.0 Build 156 04/24/2013 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_convert CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" OPERATION="INT2FLOAT" ROUNDING="TO_NEAREST" WIDTH_DATA=33 WIDTH_EXP_INPUT=8 WIDTH_EXP_OUTPUT=8 WIDTH_INT=33 WIDTH_MAN_INPUT=23 WIDTH_MAN_OUTPUT=23 WIDTH_RESULT=32 clock dataa result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:04:24:18:05:29:SJ cbx_altfp_convert 2013:04:24:18:05:29:SJ cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_altsyncram 2013:04:24:18:05:29:SJ cbx_cycloneii 2013:04:24:18:05:30:SJ cbx_lpm_abs 2013:04:24:18:05:30:SJ cbx_lpm_add_sub 2013:04:24:18:05:30:SJ cbx_lpm_compare 2013:04:24:18:05:30:SJ cbx_lpm_decode 2013:04:24:18:05:30:SJ cbx_lpm_divide 2013:04:24:18:05:30:SJ cbx_lpm_mux 2013:04:24:18:05:30:SJ cbx_mgl 2013:04:24:18:40:34:SJ cbx_stratix 2013:04:24:18:05:30:SJ cbx_stratixii 2013:04:24:18:05:30:SJ cbx_stratixiii 2013:04:24:18:05:30:SJ cbx_stratixv 2013:04:24:18:05:30:SJ cbx_util_mgl 2013:04:24:18:05:30:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" PIPELINE=2 SHIFTDIR="LEFT" SHIFTTYPE="LOGICAL" WIDTH=33 WIDTHDIST=6 aclr clk_en clock data distance result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END

--synthesis_resources = reg 71 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altbarrel_shift_drf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (32 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (32 DOWNTO 0)
	 ); 
 END altfp_convert_INT_TO_FP_altbarrel_shift_drf;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altbarrel_shift_drf IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(32 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper2d	:	STD_LOGIC_VECTOR(32 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec3r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec4r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec5r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w101w102w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w96w97w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range110w122w123w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range110w117w118w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range132w144w145w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range132w139w140w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range155w166w167w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range155w161w162w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range174w185w186w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range174w180w181w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range195w206w207w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range195w201w202w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w91w92w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range110w112w113w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range132w134w135w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range155w156w157w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range174w175w176w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range195w196w197w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range89w101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range89w96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range110w122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range110w117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range132w144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range132w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range155w166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range155w161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range174w185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range174w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range195w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range195w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range86w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range108w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range129w143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range153w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range172w184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range192w205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range89w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range110w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range132w134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range155w156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range174w175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range195w196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range89w101w102w103w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range110w122w123w124w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range132w144w145w146w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range155w166w167w168w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range174w185w186w187w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range195w206w207w208w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w104w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w125w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w147w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w169w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w188w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w209w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (230 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (197 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w116w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w120w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w138w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w142w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w160w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w164w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w179w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w183w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w200w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w204w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_pad_w_range93w_w_w_sbit_w_range84w_range94w95w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_w_sbit_w_range84w_range98w_w_pad_w_range93w99w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range149w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range171w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range190w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range84w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range107w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range127w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_smux_w_range210w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_smux_w_range148w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w101w102w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range89w101w(0) AND wire_altbarrel_shift5_w_w_w_sbit_w_range84w_range98w_w_pad_w_range93w99w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w96w97w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range89w96w(0) AND wire_altbarrel_shift5_w_w_pad_w_range93w_w_w_sbit_w_range84w_range94w95w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range110w122w123w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range110w122w(0) AND wire_altbarrel_shift5_w120w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range110w117w118w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range110w117w(0) AND wire_altbarrel_shift5_w116w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range132w144w145w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range132w144w(0) AND wire_altbarrel_shift5_w142w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range132w139w140w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range132w139w(0) AND wire_altbarrel_shift5_w138w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range155w166w167w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range155w166w(0) AND wire_altbarrel_shift5_w164w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range155w161w162w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range155w161w(0) AND wire_altbarrel_shift5_w160w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range174w185w186w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range174w185w(0) AND wire_altbarrel_shift5_w183w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range174w180w181w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range174w180w(0) AND wire_altbarrel_shift5_w179w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range195w206w207w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range195w206w(0) AND wire_altbarrel_shift5_w204w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range195w201w202w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range195w201w(0) AND wire_altbarrel_shift5_w200w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w91w92w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range89w91w(0) AND wire_altbarrel_shift5_w_sbit_w_range84w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range110w112w113w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range110w112w(0) AND wire_altbarrel_shift5_w_sbit_w_range107w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range132w134w135w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range132w134w(0) AND wire_altbarrel_shift5_w_sbit_w_range127w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range155w156w157w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range155w156w(0) AND wire_altbarrel_shift5_w_sbit_w_range149w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range174w175w176w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range174w175w(0) AND wire_altbarrel_shift5_w_sbit_w_range171w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range195w196w197w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range195w196w(0) AND wire_altbarrel_shift5_w_sbit_w_range190w(i);
	END GENERATE loop17;
	wire_altbarrel_shift5_w_lg_w_sel_w_range89w101w(0) <= wire_altbarrel_shift5_w_sel_w_range89w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range86w100w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range89w96w(0) <= wire_altbarrel_shift5_w_sel_w_range89w(0) AND wire_altbarrel_shift5_w_dir_w_range86w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range110w122w(0) <= wire_altbarrel_shift5_w_sel_w_range110w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range108w121w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range110w117w(0) <= wire_altbarrel_shift5_w_sel_w_range110w(0) AND wire_altbarrel_shift5_w_dir_w_range108w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range132w144w(0) <= wire_altbarrel_shift5_w_sel_w_range132w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range129w143w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range132w139w(0) <= wire_altbarrel_shift5_w_sel_w_range132w(0) AND wire_altbarrel_shift5_w_dir_w_range129w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range155w166w(0) <= wire_altbarrel_shift5_w_sel_w_range155w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range153w165w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range155w161w(0) <= wire_altbarrel_shift5_w_sel_w_range155w(0) AND wire_altbarrel_shift5_w_dir_w_range153w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range174w185w(0) <= wire_altbarrel_shift5_w_sel_w_range174w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range172w184w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range174w180w(0) <= wire_altbarrel_shift5_w_sel_w_range174w(0) AND wire_altbarrel_shift5_w_dir_w_range172w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range195w206w(0) <= wire_altbarrel_shift5_w_sel_w_range195w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range192w205w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range195w201w(0) <= wire_altbarrel_shift5_w_sel_w_range195w(0) AND wire_altbarrel_shift5_w_dir_w_range192w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range86w100w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range86w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range108w121w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range108w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range129w143w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range129w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range153w165w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range153w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range172w184w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range172w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range192w205w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range192w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range89w91w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range89w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range110w112w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range110w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range132w134w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range132w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range155w156w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range155w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range174w175w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range174w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range195w196w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range195w(0);
	loop18 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range89w101w102w103w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w101w102w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w96w97w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range110w122w123w124w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range110w122w123w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range110w117w118w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range132w144w145w146w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range132w144w145w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range132w139w140w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range155w166w167w168w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range155w166w167w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range155w161w162w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range174w185w186w187w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range174w185w186w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range174w180w181w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range195w206w207w208w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range195w206w207w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range195w201w202w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w104w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range89w101w102w103w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w91w92w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w125w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range110w122w123w124w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range110w112w113w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w147w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range132w144w145w146w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range132w134w135w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w169w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range155w166w167w168w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range155w156w157w(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w188w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range174w185w186w187w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range174w175w176w(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 32 GENERATE 
		wire_altbarrel_shift5_w209w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range195w206w207w208w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range195w196w197w(i);
	END GENERATE loop29;
	dir_w <= ( dir_pipe(1) & dir_w(4 DOWNTO 3) & dir_pipe(0) & dir_w(1 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(230 DOWNTO 198);
	sbit_w <= ( sbit_piper2d & smux_w(164 DOWNTO 99) & sbit_piper1d & smux_w(65 DOWNTO 0) & data);
	sel_w <= ( sel_pipec5r1d & sel_pipec4r1d & sel_pipec3r1d & distance(2 DOWNTO 0));
	smux_w <= ( wire_altbarrel_shift5_w209w & wire_altbarrel_shift5_w188w & wire_altbarrel_shift5_w169w & wire_altbarrel_shift5_w147w & wire_altbarrel_shift5_w125w & wire_altbarrel_shift5_w104w);
	wire_altbarrel_shift5_w116w <= ( pad_w(1 DOWNTO 0) & sbit_w(65 DOWNTO 35));
	wire_altbarrel_shift5_w120w <= ( sbit_w(63 DOWNTO 33) & pad_w(1 DOWNTO 0));
	wire_altbarrel_shift5_w138w <= ( pad_w(3 DOWNTO 0) & sbit_w(98 DOWNTO 70));
	wire_altbarrel_shift5_w142w <= ( sbit_w(94 DOWNTO 66) & pad_w(3 DOWNTO 0));
	wire_altbarrel_shift5_w160w <= ( pad_w(7 DOWNTO 0) & sbit_w(131 DOWNTO 107));
	wire_altbarrel_shift5_w164w <= ( sbit_w(123 DOWNTO 99) & pad_w(7 DOWNTO 0));
	wire_altbarrel_shift5_w179w <= ( pad_w(15 DOWNTO 0) & sbit_w(164 DOWNTO 148));
	wire_altbarrel_shift5_w183w <= ( sbit_w(148 DOWNTO 132) & pad_w(15 DOWNTO 0));
	wire_altbarrel_shift5_w200w <= ( pad_w(31 DOWNTO 0) & sbit_w(197));
	wire_altbarrel_shift5_w204w <= ( sbit_w(165) & pad_w(31 DOWNTO 0));
	wire_altbarrel_shift5_w_w_pad_w_range93w_w_w_sbit_w_range84w_range94w95w <= ( pad_w(0) & sbit_w(32 DOWNTO 1));
	wire_altbarrel_shift5_w_w_w_sbit_w_range84w_range98w_w_pad_w_range93w99w <= ( sbit_w(31 DOWNTO 0) & pad_w(0));
	wire_altbarrel_shift5_w_dir_w_range86w(0) <= dir_w(0);
	wire_altbarrel_shift5_w_dir_w_range108w(0) <= dir_w(1);
	wire_altbarrel_shift5_w_dir_w_range129w(0) <= dir_w(2);
	wire_altbarrel_shift5_w_dir_w_range153w(0) <= dir_w(3);
	wire_altbarrel_shift5_w_dir_w_range172w(0) <= dir_w(4);
	wire_altbarrel_shift5_w_dir_w_range192w(0) <= dir_w(5);
	wire_altbarrel_shift5_w_sbit_w_range149w <= sbit_w(131 DOWNTO 99);
	wire_altbarrel_shift5_w_sbit_w_range171w <= sbit_w(164 DOWNTO 132);
	wire_altbarrel_shift5_w_sbit_w_range190w <= sbit_w(197 DOWNTO 165);
	wire_altbarrel_shift5_w_sbit_w_range84w <= sbit_w(32 DOWNTO 0);
	wire_altbarrel_shift5_w_sbit_w_range107w <= sbit_w(65 DOWNTO 33);
	wire_altbarrel_shift5_w_sbit_w_range127w <= sbit_w(98 DOWNTO 66);
	wire_altbarrel_shift5_w_sel_w_range89w(0) <= sel_w(0);
	wire_altbarrel_shift5_w_sel_w_range110w(0) <= sel_w(1);
	wire_altbarrel_shift5_w_sel_w_range132w(0) <= sel_w(2);
	wire_altbarrel_shift5_w_sel_w_range155w(0) <= sel_w(3);
	wire_altbarrel_shift5_w_sel_w_range174w(0) <= sel_w(4);
	wire_altbarrel_shift5_w_sel_w_range195w(0) <= sel_w(5);
	wire_altbarrel_shift5_w_smux_w_range210w <= smux_w(197 DOWNTO 165);
	wire_altbarrel_shift5_w_smux_w_range148w <= smux_w(98 DOWNTO 66);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe <= ( dir_w(5) & dir_w(2));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_altbarrel_shift5_w_smux_w_range148w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper2d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper2d <= wire_altbarrel_shift5_w_smux_w_range210w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec3r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec3r1d <= distance(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec4r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec4r1d <= distance(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec5r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec5r1d <= distance(5);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --altfp_convert_INT_TO_FP_altbarrel_shift_drf


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=64 WIDTHAD=6 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END altfp_convert_INT_TO_FP_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --altfp_convert_INT_TO_FP_altpriority_encoder_3e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END altfp_convert_INT_TO_FP_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder17_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero256w257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero258w259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder18_w_lg_zero256w & wire_altpriority_encoder18_w_lg_w_lg_zero258w259w);
	zero <= (wire_altpriority_encoder17_zero AND wire_altpriority_encoder18_zero);
	altpriority_encoder17 :  altfp_convert_INT_TO_FP_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder17_q,
		zero => wire_altpriority_encoder17_zero
	  );
	wire_altpriority_encoder18_w_lg_w_lg_zero256w257w(0) <= wire_altpriority_encoder18_w_lg_zero256w(0) AND wire_altpriority_encoder18_q(0);
	wire_altpriority_encoder18_w_lg_zero258w(0) <= wire_altpriority_encoder18_zero AND wire_altpriority_encoder17_q(0);
	wire_altpriority_encoder18_w_lg_zero256w(0) <= NOT wire_altpriority_encoder18_zero;
	wire_altpriority_encoder18_w_lg_w_lg_zero258w259w(0) <= wire_altpriority_encoder18_w_lg_zero258w(0) OR wire_altpriority_encoder18_w_lg_w_lg_zero256w257w(0);
	altpriority_encoder18 :  altfp_convert_INT_TO_FP_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder18_q,
		zero => wire_altpriority_encoder18_zero
	  );

 END RTL; --altfp_convert_INT_TO_FP_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END altfp_convert_INT_TO_FP_altpriority_encoder_be8;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero246w247w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero248w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero248w249w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder16_w_lg_zero246w & wire_altpriority_encoder16_w_lg_w_lg_zero248w249w);
	zero <= (wire_altpriority_encoder15_zero AND wire_altpriority_encoder16_zero);
	altpriority_encoder15 :  altfp_convert_INT_TO_FP_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder15_q,
		zero => wire_altpriority_encoder15_zero
	  );
	loop30 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder16_w_lg_w_lg_zero246w247w(i) <= wire_altpriority_encoder16_w_lg_zero246w(0) AND wire_altpriority_encoder16_q(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder16_w_lg_zero248w(i) <= wire_altpriority_encoder16_zero AND wire_altpriority_encoder15_q(i);
	END GENERATE loop31;
	wire_altpriority_encoder16_w_lg_zero246w(0) <= NOT wire_altpriority_encoder16_zero;
	loop32 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder16_w_lg_w_lg_zero248w249w(i) <= wire_altpriority_encoder16_w_lg_zero248w(i) OR wire_altpriority_encoder16_w_lg_w_lg_zero246w247w(i);
	END GENERATE loop32;
	altpriority_encoder16 :  altfp_convert_INT_TO_FP_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder16_q,
		zero => wire_altpriority_encoder16_zero
	  );

 END RTL; --altfp_convert_INT_TO_FP_altpriority_encoder_be8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altpriority_encoder_rf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END altfp_convert_INT_TO_FP_altpriority_encoder_rf8;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altpriority_encoder_rf8 IS

	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero236w237w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero238w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero238w239w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder14_w_lg_zero236w & wire_altpriority_encoder14_w_lg_w_lg_zero238w239w);
	zero <= (wire_altpriority_encoder13_zero AND wire_altpriority_encoder14_zero);
	altpriority_encoder13 :  altfp_convert_INT_TO_FP_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );
	loop33 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero236w237w(i) <= wire_altpriority_encoder14_w_lg_zero236w(0) AND wire_altpriority_encoder14_q(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder14_w_lg_zero238w(i) <= wire_altpriority_encoder14_zero AND wire_altpriority_encoder13_q(i);
	END GENERATE loop34;
	wire_altpriority_encoder14_w_lg_zero236w(0) <= NOT wire_altpriority_encoder14_zero;
	loop35 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero238w239w(i) <= wire_altpriority_encoder14_w_lg_zero238w(i) OR wire_altpriority_encoder14_w_lg_w_lg_zero236w237w(i);
	END GENERATE loop35;
	altpriority_encoder14 :  altfp_convert_INT_TO_FP_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder14_q,
		zero => wire_altpriority_encoder14_zero
	  );

 END RTL; --altfp_convert_INT_TO_FP_altpriority_encoder_rf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altpriority_encoder_qf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END altfp_convert_INT_TO_FP_altpriority_encoder_qf8;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altpriority_encoder_qf8 IS

	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero226w227w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero228w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero228w229w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder12_w_lg_zero226w & wire_altpriority_encoder12_w_lg_w_lg_zero228w229w);
	zero <= (wire_altpriority_encoder11_zero AND wire_altpriority_encoder12_zero);
	altpriority_encoder11 :  altfp_convert_INT_TO_FP_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );
	loop36 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder12_w_lg_w_lg_zero226w227w(i) <= wire_altpriority_encoder12_w_lg_zero226w(0) AND wire_altpriority_encoder12_q(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder12_w_lg_zero228w(i) <= wire_altpriority_encoder12_zero AND wire_altpriority_encoder11_q(i);
	END GENERATE loop37;
	wire_altpriority_encoder12_w_lg_zero226w(0) <= NOT wire_altpriority_encoder12_zero;
	loop38 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder12_w_lg_w_lg_zero228w229w(i) <= wire_altpriority_encoder12_w_lg_zero228w(i) OR wire_altpriority_encoder12_w_lg_w_lg_zero226w227w(i);
	END GENERATE loop38;
	altpriority_encoder12 :  altfp_convert_INT_TO_FP_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder12_q,
		zero => wire_altpriority_encoder12_zero
	  );

 END RTL; --altfp_convert_INT_TO_FP_altpriority_encoder_qf8


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:04:24:18:05:29:SJ cbx_mgl 2013:04:24:18:40:34:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END altfp_convert_INT_TO_FP_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --altfp_convert_INT_TO_FP_altpriority_encoder_3v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END altfp_convert_INT_TO_FP_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder25_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder26_w_lg_w_lg_zero299w300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder26_w_lg_zero301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder26_w_lg_zero299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder26_w_lg_w_lg_zero301w302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder26_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder26_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder26_w_lg_zero299w & wire_altpriority_encoder26_w_lg_w_lg_zero301w302w);
	altpriority_encoder25 :  altfp_convert_INT_TO_FP_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder25_q
	  );
	wire_altpriority_encoder26_w_lg_w_lg_zero299w300w(0) <= wire_altpriority_encoder26_w_lg_zero299w(0) AND wire_altpriority_encoder26_q(0);
	wire_altpriority_encoder26_w_lg_zero301w(0) <= wire_altpriority_encoder26_zero AND wire_altpriority_encoder25_q(0);
	wire_altpriority_encoder26_w_lg_zero299w(0) <= NOT wire_altpriority_encoder26_zero;
	wire_altpriority_encoder26_w_lg_w_lg_zero301w302w(0) <= wire_altpriority_encoder26_w_lg_zero301w(0) OR wire_altpriority_encoder26_w_lg_w_lg_zero299w300w(0);
	altpriority_encoder26 :  altfp_convert_INT_TO_FP_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder26_q,
		zero => wire_altpriority_encoder26_zero
	  );

 END RTL; --altfp_convert_INT_TO_FP_altpriority_encoder_6v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END altfp_convert_INT_TO_FP_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder23_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_w_lg_w_lg_zero290w291w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_w_lg_zero292w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_w_lg_zero290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_w_lg_w_lg_zero292w293w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder24_w_lg_zero290w & wire_altpriority_encoder24_w_lg_w_lg_zero292w293w);
	altpriority_encoder23 :  altfp_convert_INT_TO_FP_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder23_q
	  );
	loop39 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder24_w_lg_w_lg_zero290w291w(i) <= wire_altpriority_encoder24_w_lg_zero290w(0) AND wire_altpriority_encoder24_q(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder24_w_lg_zero292w(i) <= wire_altpriority_encoder24_zero AND wire_altpriority_encoder23_q(i);
	END GENERATE loop40;
	wire_altpriority_encoder24_w_lg_zero290w(0) <= NOT wire_altpriority_encoder24_zero;
	loop41 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder24_w_lg_w_lg_zero292w293w(i) <= wire_altpriority_encoder24_w_lg_zero292w(i) OR wire_altpriority_encoder24_w_lg_w_lg_zero290w291w(i);
	END GENERATE loop41;
	altpriority_encoder24 :  altfp_convert_INT_TO_FP_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder24_q,
		zero => wire_altpriority_encoder24_zero
	  );

 END RTL; --altfp_convert_INT_TO_FP_altpriority_encoder_bv7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altpriority_encoder_r08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END altfp_convert_INT_TO_FP_altpriority_encoder_r08;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altpriority_encoder_r08 IS

	 SIGNAL  wire_altpriority_encoder21_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero281w282w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero283w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero283w284w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder22_w_lg_zero281w & wire_altpriority_encoder22_w_lg_w_lg_zero283w284w);
	altpriority_encoder21 :  altfp_convert_INT_TO_FP_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder21_q
	  );
	loop42 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder22_w_lg_w_lg_zero281w282w(i) <= wire_altpriority_encoder22_w_lg_zero281w(0) AND wire_altpriority_encoder22_q(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder22_w_lg_zero283w(i) <= wire_altpriority_encoder22_zero AND wire_altpriority_encoder21_q(i);
	END GENERATE loop43;
	wire_altpriority_encoder22_w_lg_zero281w(0) <= NOT wire_altpriority_encoder22_zero;
	loop44 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder22_w_lg_w_lg_zero283w284w(i) <= wire_altpriority_encoder22_w_lg_zero283w(i) OR wire_altpriority_encoder22_w_lg_w_lg_zero281w282w(i);
	END GENERATE loop44;
	altpriority_encoder22 :  altfp_convert_INT_TO_FP_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder22_q,
		zero => wire_altpriority_encoder22_zero
	  );

 END RTL; --altfp_convert_INT_TO_FP_altpriority_encoder_r08

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altpriority_encoder_q08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END altfp_convert_INT_TO_FP_altpriority_encoder_q08;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altpriority_encoder_q08 IS

	 SIGNAL  wire_altpriority_encoder19_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero272w273w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero274w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero274w275w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder20_w_lg_zero272w & wire_altpriority_encoder20_w_lg_w_lg_zero274w275w);
	altpriority_encoder19 :  altfp_convert_INT_TO_FP_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder19_q
	  );
	loop45 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero272w273w(i) <= wire_altpriority_encoder20_w_lg_zero272w(0) AND wire_altpriority_encoder20_q(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_zero274w(i) <= wire_altpriority_encoder20_zero AND wire_altpriority_encoder19_q(i);
	END GENERATE loop46;
	wire_altpriority_encoder20_w_lg_zero272w(0) <= NOT wire_altpriority_encoder20_zero;
	loop47 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero274w275w(i) <= wire_altpriority_encoder20_w_lg_zero274w(i) OR wire_altpriority_encoder20_w_lg_w_lg_zero272w273w(i);
	END GENERATE loop47;
	altpriority_encoder20 :  altfp_convert_INT_TO_FP_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder20_q,
		zero => wire_altpriority_encoder20_zero
	  );

 END RTL; --altfp_convert_INT_TO_FP_altpriority_encoder_q08

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altpriority_encoder_0c6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0)
	 ); 
 END altfp_convert_INT_TO_FP_altpriority_encoder_0c6;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altpriority_encoder_0c6 IS

	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero217w218w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero219w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero219w220w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_qf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_q08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder10_w_lg_zero217w & wire_altpriority_encoder10_w_lg_w_lg_zero219w220w);
	loop48 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder10_w_lg_w_lg_zero217w218w(i) <= wire_altpriority_encoder10_w_lg_zero217w(0) AND wire_altpriority_encoder10_q(i);
	END GENERATE loop48;
	loop49 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder10_w_lg_zero219w(i) <= wire_altpriority_encoder10_zero AND wire_altpriority_encoder9_q(i);
	END GENERATE loop49;
	wire_altpriority_encoder10_w_lg_zero217w(0) <= NOT wire_altpriority_encoder10_zero;
	loop50 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder10_w_lg_w_lg_zero219w220w(i) <= wire_altpriority_encoder10_w_lg_zero219w(i) OR wire_altpriority_encoder10_w_lg_w_lg_zero217w218w(i);
	END GENERATE loop50;
	altpriority_encoder10 :  altfp_convert_INT_TO_FP_altpriority_encoder_qf8
	  PORT MAP ( 
		data => data(63 DOWNTO 32),
		q => wire_altpriority_encoder10_q,
		zero => wire_altpriority_encoder10_zero
	  );
	altpriority_encoder9 :  altfp_convert_INT_TO_FP_altpriority_encoder_q08
	  PORT MAP ( 
		data => data(31 DOWNTO 0),
		q => wire_altpriority_encoder9_q
	  );

 END RTL; --altfp_convert_INT_TO_FP_altpriority_encoder_0c6

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 5 lpm_compare 1 reg 253 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert_INT_TO_FP_altfp_convert_5tm IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (32 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END altfp_convert_INT_TO_FP_altfp_convert_5tm;

 ARCHITECTURE RTL OF altfp_convert_INT_TO_FP_altfp_convert_5tm IS

	 SIGNAL  wire_altbarrel_shift5_data	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_result	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder2_data	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder2_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL	 add_1_adder1_cout_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_w_lg_q64w65w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_q62w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_q64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 add_1_adder1_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_adder2_cout_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_adder2_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_1_reg_w_lg_w_lg_q71w72w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_1_reg_w_lg_q70w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_1_reg_w_lg_q71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exponent_bus_pre_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg2	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissa_pre_round_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_mantissa_pre_round_reg_w_q_range63w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL	 priority_encoder_reg	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 result_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub1_datab	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub6_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub6_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub6_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub7_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub7_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub7_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub8_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub8_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_w_lg_alb22w23w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_alb21w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_alb22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cmpr4_alb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_guard_bit_w56w57w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_guard_bit_w56w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mantissa_overflow75w76w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_max_neg_value_selector18w19w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_int_a5w6w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_mantissa_overflow74w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector17w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a4w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_guard_bit_w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mantissa_overflow75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range35w38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range39w41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range42w44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range45w47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range48w50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range51w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  add_1_adder1_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  add_1_adder2_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  add_1_adder_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  add_1_w :	STD_LOGIC;
	 SIGNAL  bias_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  const_bias_value_add_width_int_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exceptions_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_bus :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_bus_pre :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_output_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_rounded :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  guard_bit_w :	STD_LOGIC;
	 SIGNAL  int_a :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  int_a_2s :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  invert_int_a :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  leading_zeroes :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  mag_int_a :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  mantissa_bus :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  mantissa_overflow :	STD_LOGIC;
	 SIGNAL  mantissa_post_round :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  mantissa_pre_round :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  mantissa_rounded :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  max_neg_value_selector :	STD_LOGIC;
	 SIGNAL  max_neg_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  minus_leading_zero :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  prio_mag_int_a :	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  priority_pad_one_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  round_bit_w :	STD_LOGIC;
	 SIGNAL  shifted_mag_int_a :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  sign_bus :	STD_LOGIC;
	 SIGNAL  sign_int_a :	STD_LOGIC;
	 SIGNAL  sticky_bit_bus :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  sticky_bit_or_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  sticky_bit_w :	STD_LOGIC;
	 SIGNAL  zero_padding_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  altfp_convert_INT_TO_FP_altbarrel_shift_drf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(32 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(32 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altfp_convert_INT_TO_FP_altpriority_encoder_0c6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_guard_bit_w56w57w58w(0) <= wire_w_lg_w_lg_guard_bit_w56w57w(0) AND sticky_bit_w;
	wire_w_lg_w_lg_guard_bit_w56w57w(0) <= wire_w_lg_guard_bit_w56w(0) AND round_bit_w;
	loop51 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_mantissa_overflow75w76w(i) <= wire_w_lg_mantissa_overflow75w(0) AND exponent_bus_pre_reg(i);
	END GENERATE loop51;
	loop52 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_max_neg_value_selector18w19w(i) <= wire_w_lg_max_neg_value_selector18w(0) AND exponent_zero_w(i);
	END GENERATE loop52;
	loop53 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_lg_sign_int_a5w6w(i) <= wire_w_lg_sign_int_a5w(0) AND int_a(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_mantissa_overflow74w(i) <= mantissa_overflow AND wire_add_sub8_result(i);
	END GENERATE loop54;
	loop55 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_max_neg_value_selector17w(i) <= max_neg_value_selector AND max_neg_value_w(i);
	END GENERATE loop55;
	loop56 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_sign_int_a4w(i) <= sign_int_a AND int_a_2s(i);
	END GENERATE loop56;
	wire_w_lg_guard_bit_w56w(0) <= NOT guard_bit_w;
	wire_w_lg_mantissa_overflow75w(0) <= NOT mantissa_overflow;
	wire_w_lg_max_neg_value_selector18w(0) <= NOT max_neg_value_selector;
	wire_w_lg_sign_int_a5w(0) <= NOT sign_int_a;
	wire_w_lg_w_sticky_bit_or_w_range35w38w(0) <= wire_w_sticky_bit_or_w_range35w(0) OR wire_w_sticky_bit_bus_range37w(0);
	wire_w_lg_w_sticky_bit_or_w_range39w41w(0) <= wire_w_sticky_bit_or_w_range39w(0) OR wire_w_sticky_bit_bus_range40w(0);
	wire_w_lg_w_sticky_bit_or_w_range42w44w(0) <= wire_w_sticky_bit_or_w_range42w(0) OR wire_w_sticky_bit_bus_range43w(0);
	wire_w_lg_w_sticky_bit_or_w_range45w47w(0) <= wire_w_sticky_bit_or_w_range45w(0) OR wire_w_sticky_bit_bus_range46w(0);
	wire_w_lg_w_sticky_bit_or_w_range48w50w(0) <= wire_w_sticky_bit_or_w_range48w(0) OR wire_w_sticky_bit_bus_range49w(0);
	wire_w_lg_w_sticky_bit_or_w_range51w53w(0) <= wire_w_sticky_bit_or_w_range51w(0) OR wire_w_sticky_bit_bus_range52w(0);
	aclr <= '0';
	add_1_adder1_w <= add_1_adder1_reg;
	add_1_adder2_w <= (wire_add_1_adder1_cout_reg_w_lg_w_lg_q64w65w OR wire_add_1_adder1_cout_reg_w_lg_q62w);
	add_1_adder_w <= ( add_1_adder2_w & add_1_adder1_w);
	add_1_w <= (wire_w_lg_w_lg_w_lg_guard_bit_w56w57w58w(0) OR (guard_bit_w AND round_bit_w));
	bias_value_w <= "01111111";
	clk_en <= '1';
	const_bias_value_add_width_int_w <= "10011110";
	exceptions_value <= (wire_w_lg_w_lg_max_neg_value_selector18w19w OR wire_w_lg_max_neg_value_selector17w);
	exponent_bus <= exponent_rounded;
	exponent_bus_pre <= (wire_cmpr4_w_lg_w_lg_alb22w23w OR wire_cmpr4_w_lg_alb21w);
	exponent_output_w <= wire_add_sub3_result;
	exponent_rounded <= (wire_w_lg_w_lg_mantissa_overflow75w76w OR wire_w_lg_mantissa_overflow74w);
	exponent_zero_w <= (OTHERS => '0');
	guard_bit_w <= shifted_mag_int_a(8);
	int_a <= dataa(31 DOWNTO 0);
	int_a_2s <= wire_add_sub1_result;
	invert_int_a <= (NOT int_a);
	leading_zeroes <= (NOT priority_encoder_reg);
	mag_int_a <= (wire_w_lg_w_lg_sign_int_a5w6w OR wire_w_lg_sign_int_a4w);
	mantissa_bus <= mantissa_rounded(22 DOWNTO 0);
	mantissa_overflow <= ((add_1_reg AND add_1_adder1_cout_reg) AND add_1_adder2_cout_reg);
	mantissa_post_round <= add_1_adder_w;
	mantissa_pre_round <= shifted_mag_int_a(31 DOWNTO 8);
	mantissa_rounded <= (wire_add_1_reg_w_lg_w_lg_q71w72w OR wire_add_1_reg_w_lg_q70w);
	max_neg_value_selector <= (wire_cmpr4_alb AND sign_int_a_reg2);
	max_neg_value_w <= "10011111";
	minus_leading_zero <= ( zero_padding_w & leading_zeroes);
	prio_mag_int_a <= ( mag_int_a_reg & "1");
	priority_pad_one_w <= (OTHERS => '1');
	result <= result_reg;
	result_w <= ( sign_bus & exponent_bus & mantissa_bus);
	round_bit_w <= shifted_mag_int_a(7);
	shifted_mag_int_a <= wire_altbarrel_shift5_result(31 DOWNTO 0);
	sign_bus <= sign_int_a_reg5;
	sign_int_a <= dataa(32);
	sticky_bit_bus <= shifted_mag_int_a(6 DOWNTO 0);
	sticky_bit_or_w <= ( wire_w_lg_w_sticky_bit_or_w_range51w53w & wire_w_lg_w_sticky_bit_or_w_range48w50w & wire_w_lg_w_sticky_bit_or_w_range45w47w & wire_w_lg_w_sticky_bit_or_w_range42w44w & wire_w_lg_w_sticky_bit_or_w_range39w41w & wire_w_lg_w_sticky_bit_or_w_range35w38w & sticky_bit_bus(0));
	sticky_bit_w <= sticky_bit_or_w(6);
	zero_padding_w <= (OTHERS => '0');
	wire_w_sticky_bit_bus_range37w(0) <= sticky_bit_bus(1);
	wire_w_sticky_bit_bus_range40w(0) <= sticky_bit_bus(2);
	wire_w_sticky_bit_bus_range43w(0) <= sticky_bit_bus(3);
	wire_w_sticky_bit_bus_range46w(0) <= sticky_bit_bus(4);
	wire_w_sticky_bit_bus_range49w(0) <= sticky_bit_bus(5);
	wire_w_sticky_bit_bus_range52w(0) <= sticky_bit_bus(6);
	wire_w_sticky_bit_or_w_range35w(0) <= sticky_bit_or_w(0);
	wire_w_sticky_bit_or_w_range39w(0) <= sticky_bit_or_w(1);
	wire_w_sticky_bit_or_w_range42w(0) <= sticky_bit_or_w(2);
	wire_w_sticky_bit_or_w_range45w(0) <= sticky_bit_or_w(3);
	wire_w_sticky_bit_or_w_range48w(0) <= sticky_bit_or_w(4);
	wire_w_sticky_bit_or_w_range51w(0) <= sticky_bit_or_w(5);
	wire_altbarrel_shift5_data <= ( "0" & mag_int_a_reg2);
	altbarrel_shift5 :  altfp_convert_INT_TO_FP_altbarrel_shift_drf
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_altbarrel_shift5_data,
		distance => leading_zeroes,
		result => wire_altbarrel_shift5_result
	  );
	wire_altpriority_encoder2_data <= ( prio_mag_int_a & priority_pad_one_w);
	altpriority_encoder2 :  altfp_convert_INT_TO_FP_altpriority_encoder_0c6
	  PORT MAP ( 
		data => wire_altpriority_encoder2_data,
		q => wire_altpriority_encoder2_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder1_cout_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder1_cout_reg <= wire_add_sub6_cout;
			END IF;
		END IF;
	END PROCESS;
	loop57 : FOR i IN 0 TO 11 GENERATE 
		wire_add_1_adder1_cout_reg_w_lg_w_lg_q64w65w(i) <= wire_add_1_adder1_cout_reg_w_lg_q64w(0) AND wire_mantissa_pre_round_reg_w_q_range63w(i);
	END GENERATE loop57;
	loop58 : FOR i IN 0 TO 11 GENERATE 
		wire_add_1_adder1_cout_reg_w_lg_q62w(i) <= add_1_adder1_cout_reg AND add_1_adder2_reg(i);
	END GENERATE loop58;
	wire_add_1_adder1_cout_reg_w_lg_q64w(0) <= NOT add_1_adder1_cout_reg;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder1_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder1_reg <= wire_add_sub6_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder2_cout_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder2_cout_reg <= wire_add_sub7_cout;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder2_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder2_reg <= wire_add_sub7_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_reg <= add_1_w;
			END IF;
		END IF;
	END PROCESS;
	loop59 : FOR i IN 0 TO 23 GENERATE 
		wire_add_1_reg_w_lg_w_lg_q71w72w(i) <= wire_add_1_reg_w_lg_q71w(0) AND mantissa_pre_round_reg(i);
	END GENERATE loop59;
	loop60 : FOR i IN 0 TO 23 GENERATE 
		wire_add_1_reg_w_lg_q70w(i) <= add_1_reg AND mantissa_post_round(i);
	END GENERATE loop60;
	wire_add_1_reg_w_lg_q71w(0) <= NOT add_1_reg;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg <= exponent_bus_pre_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg2 <= exponent_bus_pre_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg3 <= exponent_bus_pre;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg <= mag_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg2 <= mag_int_a_reg;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissa_pre_round_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissa_pre_round_reg <= mantissa_pre_round;
			END IF;
		END IF;
	END PROCESS;
	wire_mantissa_pre_round_reg_w_q_range63w <= mantissa_pre_round_reg(23 DOWNTO 12);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN priority_encoder_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN priority_encoder_reg <= wire_altpriority_encoder2_q;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN result_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN result_reg <= result_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg1 <= sign_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg2 <= sign_int_a_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg3 <= sign_int_a_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg4 <= sign_int_a_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg5 <= sign_int_a_reg4;
			END IF;
		END IF;
	END PROCESS;
	wire_add_sub1_datab <= "00000000000000000000000000000001";
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 32,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => invert_int_a,
		datab => wire_add_sub1_datab,
		result => wire_add_sub1_result
	  );
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => const_bias_value_add_width_int_w,
		datab => minus_leading_zero,
		result => wire_add_sub3_result
	  );
	wire_add_sub6_datab <= "000000000001";
	add_sub6 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 12,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub6_cout,
		dataa => mantissa_pre_round(11 DOWNTO 0),
		datab => wire_add_sub6_datab,
		result => wire_add_sub6_result
	  );
	wire_add_sub7_datab <= "000000000001";
	add_sub7 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 12,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub7_cout,
		dataa => mantissa_pre_round(23 DOWNTO 12),
		datab => wire_add_sub7_datab,
		result => wire_add_sub7_result
	  );
	wire_add_sub8_datab <= "00000001";
	add_sub8 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => exponent_bus_pre_reg,
		datab => wire_add_sub8_datab,
		result => wire_add_sub8_result
	  );
	loop61 : FOR i IN 0 TO 7 GENERATE 
		wire_cmpr4_w_lg_w_lg_alb22w23w(i) <= wire_cmpr4_w_lg_alb22w(0) AND exponent_output_w(i);
	END GENERATE loop61;
	loop62 : FOR i IN 0 TO 7 GENERATE 
		wire_cmpr4_w_lg_alb21w(i) <= wire_cmpr4_alb AND exceptions_value(i);
	END GENERATE loop62;
	wire_cmpr4_w_lg_alb22w(0) <= NOT wire_cmpr4_alb;
	cmpr4 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		alb => wire_cmpr4_alb,
		dataa => exponent_output_w,
		datab => bias_value_w
	  );

 END RTL; --altfp_convert_INT_TO_FP_altfp_convert_5tm
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altfp_convert_INT_TO_FP IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (32 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END altfp_convert_INT_TO_FP;


ARCHITECTURE RTL OF altfp_convert_int_to_fp IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT altfp_convert_INT_TO_FP_altfp_convert_5tm
	PORT (
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (32 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	altfp_convert_INT_TO_FP_altfp_convert_5tm_component : altfp_convert_INT_TO_FP_altfp_convert_5tm
	PORT MAP (
		clock => clock,
		dataa => dataa,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_convert"
-- Retrieval info: CONSTANT: OPERATION STRING "INT2FLOAT"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "33"
-- Retrieval info: CONSTANT: WIDTH_EXP_INPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_EXP_OUTPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_INT NUMERIC "33"
-- Retrieval info: CONSTANT: WIDTH_MAN_INPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_MAN_OUTPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "32"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 33 0 INPUT NODEFVAL "dataa[32..0]"
-- Retrieval info: CONNECT: @dataa 0 0 33 0 dataa 0 0 33 0
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert_INT_TO_FP.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert_INT_TO_FP.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert_INT_TO_FP.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert_INT_TO_FP_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert_INT_TO_FP.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert_INT_TO_FP.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: lpm
