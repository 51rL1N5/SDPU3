altfp_convert_INT_TO_FP_inst : altfp_convert_INT_TO_FP PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
