library verilog;
use verilog.vl_types.all;
entity Secador_vlg_vec_tst is
end Secador_vlg_vec_tst;
