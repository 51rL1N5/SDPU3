altfp_mult_ADJUSTING_DATA_inst : altfp_mult_ADJUSTING_DATA PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
