altfp_convert_FP_TO_INT_inst : altfp_convert_FP_TO_INT PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
